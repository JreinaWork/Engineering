*Vacuum Tube Triode (Audio freq.) pkg:VT-9 (A:1,2,3)(B:6,7,8)
*Connections:
*             Plate
*             | Grid
*             | | Cathode
*             | | |
.SUBCKT 12AX7 1 3 4
B1 2 4 I=((URAMP((V(2,4)/85)+V(3,4)))^1.5)/580
C1 3 4 1.6E-12
C2 3 1 1.7E-12
C3 1 4 0.46E-12
R1 3 5 50E+3
D1 1 2 DX
D2 4 2 DX2
D3 5 4 DX
.MODEL DX D(IS=1.0E-12 RS=1.0)
.MODEL DX2 D(IS=1.0E-9 RS=1.0)
.ENDS X12AX7

*LF411C
*Sngl LoOffset LoDrift JFET OpAmp pkg:DIP8 3,2,8,4,6. pkg:CAN8 3,2,8,4,6.
*
* Connections:
*               Non-Inverting Input
*               | Inverting Input
*               | | Positive Power Supply
*               | | | Negative Power Supply
*               | | | | Output
*               | | | | |
.SUBCKT LF411C  1 2 3 4 5
  C1   11 12 3.498E-12
  C2    6  7 15E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  BGND 99  0 V=V(3)*.5 + V(4)*.5
  BB    7 99 I=I(VB)*28.29E6 - I(VC)*30E6 + I(VE)*30E6 +
+              I(VLP)*30E6 - I(VLN)*30E6
  GA    6  0 11 12 282.8E-6
  GCM   0  6 10 99 1.59E-9
  ISS   3 10 DC 195E-6
  HLIM 90  0 VLIM 1K
  J1   11  2 10 JX
  J2   12  1 10 JX
  R2    6  9 100E3
  RD1   4 11 3.536E3
  RD2   4 12 3.536E3
  RO1   8  5 50
  RO2   7 99 25
  RP    3  4 15E3
  RSS  10 99 1.026E6
  VB    9  0 DC 0
  VC    3 53 DC 2.2
  VE   54  4 DC 2.2
  VLIM  7  8 DC 0
  VLP  91  0 DC 30
  VLN   0 92 DC 30
.MODEL DX D(IS=800E-18)
.MODEL JX PJF(IS=12.5E-12 BETA=250.1E-6 VTO=-1)
.ENDS LF411C
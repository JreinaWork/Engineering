*Crystal Subcircuit Parameters
*FREQ = Fundamental frequency 
*RS   = Series resistance
*C    = Parallel capacitance
*Q    = Quality Factor

*CTS Color Burst alias:XCRYSTAL {FREQ=3.58E6 RS=160 C=1.8E-11} pkg:HC49	
.SUBCKT 3.5795MHZ 1 2 PARAMS: FREQ=3.58E6 RS=160 C=1.8E-11 Q=1000
LX 1 3 {((Q*RS)/(6.2831852*FREQ))} IC=0.5M
CX 3 4 {(1/(Q*6.2831852*FREQ*RS))}
C0 1 2 {C}
RS 4 2 {RS}
.ENDS

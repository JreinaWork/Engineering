*====================================================
*uA741
*Sngl GenPurpose OpAmp pkg:DIP8 3,2,7,4,6. pkg:CAN8 3,2,7,4,6.
* Connections: 
*             Non-Inverting Input
*             | Inverting Input
*             | | Positive Power Supply
*             | | | Negative Power Supply
*             | | | | Output
*             | | | | |
.SUBCKT UA741 1 2 3 4 5
  C1   11 12 4.664E-12
  C2    6  7 20E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  BGND 99  0 V=V(3)*.5 + V(4)*.5
  BB    7 99 I=I(VB)*10.61E6 - I(VC)*10E6 + I(VE)*10E6 +
+              I(VLP)*10E6 - I(VLN)*10E6
  GA    6  0 11 12 137.7E-6
  GCM   0  6 10 99 2.574E-9
  IEE  10  4 DC 10.16E-6
  HLIM 90  0 VLIM 1K
  Q1   11  2 13 QX
  Q2   12  1 14 QX
  R2    6  9 100E3
  RC1   3 11 7.957E3
  RC2   3 12 7.957E3
  RE1  13 10 2.74E3
  RE2  14 10 2.74E3
  REE  10 99 19.69E6
  RO1   8  5 150
  RO2   7 99 150
  RP    3  4 18.11E3
  VB    9  0 DC 0
  VC    3 53 DC 2.6
  VE   54  4 DC 2.6
  VLIM  7  8 DC 0
  VLP  91  0 DC 25
  VLN   0 92 DC 25
.MODEL DX D(IS=800E-18)
.MODEL QX NPN(IS=800E-18 BF=62.5)
.ENDS UA741

* Origin: Mcemods2.lib

*18DB10 MCE 4-8-96
*Ref: IR Power Semiconductors Product Digest '94
*1000V 1.8A Si pkg:D-2
.SUBCKT 18DB10 1 2 3 4
D1 1 2 18DB10
D2 1 4 18DB10
D3 2 3 18DB10
D4 4 3 18DB10
.MODEL 18DB10 D (IS=4.94N RS=42M N=1.75 BV=1K IBV=191U
+ CJO=75.3P VJ=.75 M=.333 TT=4.32U)
.ENDS D18DB10

* Origin: Mcediode.lib
